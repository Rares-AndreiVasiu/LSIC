module display7bit(
	input [3 : 0] cnt,
	output [ 7 : 0]
